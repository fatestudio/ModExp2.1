`include "_parameter.v"

module ModExp_tb();
	reg clk;
	reg reset;
	reg [`DATA_WIDTH16 - 1 : 0] m_buf;
	reg [`DATA_WIDTH16 - 1 : 0] e_buf;
	reg [`DATA_WIDTH16 - 1 : 0] n_buf;
	reg [`DATA_WIDTH16 - 1 : 0] r_buf;
	reg [`DATA_WIDTH16 - 1 : 0] t_buf;
	reg [`DATA_WIDTH16 - 1 : 0] nprime0_buf;
	reg startInput;
	reg startCompute;
	reg getResult;
	wire [`DATA_WIDTH16 - 1 : 0] res_out;
	wire [4 : 0] exp_state;
	wire [3 : 0] state;
	
	ModExp modexp0(
		.clk(clk), .reset(reset), .m_buf(m_buf), .e_buf(e_buf), .n_buf(n_buf), .r_buf(r_buf), .t_buf(t_buf), .nprime0_buf(nprime0_buf),
		.startInput(startInput), .startCompute(startCompute), .getResult(getResult), 
		.exp_state(exp_state), .state(state), .res_out(res_out)
	);
	
	initial begin
		clk = 0;
		reset = 0;
		startInput = 0;
		startCompute = 0;
		getResult = 0;
		m_buf = 16'h0000;
		e_buf = 16'h0000;
		n_buf = 16'h0000;
		r_buf = 16'h0000;
		t_buf = 16'h0000;
		nprime0_buf = 16'h0000;
		#100 
		startInput = 1;	

#10
m_buf = 16'h6d1d;
e_buf = 16'h0005;
n_buf = 16'h898f;
r_buf = 16'h7671;
t_buf = 16'h289e;
nprime0_buf = 16'h8a91;
#10
m_buf = 16'h42cb;
e_buf = 16'h0000;
n_buf = 16'h5fec;
r_buf = 16'ha013;
t_buf = 16'hacaa;
nprime0_buf = 16'ha3b1;
#10
m_buf = 16'h8051;
e_buf = 16'h0000;
n_buf = 16'hbd79;
r_buf = 16'h4286;
t_buf = 16'h3f82;
nprime0_buf = 16'h2df6;
#10
m_buf = 16'h95d1;
e_buf = 16'h0000;
n_buf = 16'h1622;
r_buf = 16'he9dd;
t_buf = 16'h7305;
nprime0_buf = 16'h3bea;
#10
m_buf = 16'h0933;
e_buf = 16'h0000;
n_buf = 16'hca16;
r_buf = 16'h35e9;
t_buf = 16'hf2c5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc6f0;
e_buf = 16'h0000;
n_buf = 16'h705f;
r_buf = 16'h8fa0;
t_buf = 16'h2b90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0f4e;
e_buf = 16'h0000;
n_buf = 16'h0806;
r_buf = 16'hf7f9;
t_buf = 16'h6657;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2aa5;
e_buf = 16'h0000;
n_buf = 16'ha9ec;
r_buf = 16'h5613;
t_buf = 16'h4906;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8043;
e_buf = 16'h0000;
n_buf = 16'h3d15;
r_buf = 16'hc2ea;
t_buf = 16'h0a06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6e64;
e_buf = 16'h0000;
n_buf = 16'h8228;
r_buf = 16'h7dd7;
t_buf = 16'h0040;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4efe;
e_buf = 16'h0000;
n_buf = 16'h6215;
r_buf = 16'h9dea;
t_buf = 16'h0115;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3123;
e_buf = 16'h0000;
n_buf = 16'h1ba1;
r_buf = 16'he45e;
t_buf = 16'h41d7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfdeb;
e_buf = 16'h0000;
n_buf = 16'h03e3;
r_buf = 16'hfc1c;
t_buf = 16'h4bdb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5bc7;
e_buf = 16'h0000;
n_buf = 16'hc748;
r_buf = 16'h38b7;
t_buf = 16'hd1a3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h73e5;
e_buf = 16'h0000;
n_buf = 16'h21a4;
r_buf = 16'hde5b;
t_buf = 16'hb841;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1d71;
e_buf = 16'h0000;
n_buf = 16'h29e8;
r_buf = 16'hd617;
t_buf = 16'h4255;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfe8c;
e_buf = 16'h0000;
n_buf = 16'h3844;
r_buf = 16'hc7bb;
t_buf = 16'h73e0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1058;
e_buf = 16'h0000;
n_buf = 16'h855c;
r_buf = 16'h7aa3;
t_buf = 16'hdf44;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5396;
e_buf = 16'h0000;
n_buf = 16'h107e;
r_buf = 16'hef81;
t_buf = 16'hbcdf;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd26d;
e_buf = 16'h0000;
n_buf = 16'hd707;
r_buf = 16'h28f8;
t_buf = 16'h0d21;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8266;
e_buf = 16'h0000;
n_buf = 16'h5db9;
r_buf = 16'ha246;
t_buf = 16'hfa55;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdd13;
e_buf = 16'h0000;
n_buf = 16'h64ac;
r_buf = 16'h9b53;
t_buf = 16'h386e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf267;
e_buf = 16'h0000;
n_buf = 16'h92d8;
r_buf = 16'h6d27;
t_buf = 16'hce5f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hda54;
e_buf = 16'h0000;
n_buf = 16'h5eda;
r_buf = 16'ha125;
t_buf = 16'hef79;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8b57;
e_buf = 16'h0000;
n_buf = 16'h8dfc;
r_buf = 16'h7203;
t_buf = 16'h8c2e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3b6;
e_buf = 16'h0000;
n_buf = 16'h7d5c;
r_buf = 16'h82a3;
t_buf = 16'h2b88;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0911;
e_buf = 16'h0000;
n_buf = 16'h8a43;
r_buf = 16'h75bc;
t_buf = 16'hbaa2;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0712;
e_buf = 16'h0000;
n_buf = 16'hbb96;
r_buf = 16'h4469;
t_buf = 16'ha401;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb5b7;
e_buf = 16'h0000;
n_buf = 16'h3986;
r_buf = 16'hc679;
t_buf = 16'hf001;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he72b;
e_buf = 16'h0000;
n_buf = 16'h0792;
r_buf = 16'hf86d;
t_buf = 16'h0135;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdbd2;
e_buf = 16'h0000;
n_buf = 16'h5d68;
r_buf = 16'ha297;
t_buf = 16'h1e91;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h869b;
e_buf = 16'h0000;
n_buf = 16'h7825;
r_buf = 16'h87da;
t_buf = 16'h432c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd488;
e_buf = 16'h0000;
n_buf = 16'hfbac;
r_buf = 16'h0453;
t_buf = 16'hd484;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h739c;
e_buf = 16'h0000;
n_buf = 16'h0b21;
r_buf = 16'hf4de;
t_buf = 16'h9f25;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcd8f;
e_buf = 16'h0000;
n_buf = 16'hc8d6;
r_buf = 16'h3729;
t_buf = 16'h6bf1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc09f;
e_buf = 16'h0000;
n_buf = 16'h4efb;
r_buf = 16'hb104;
t_buf = 16'h192d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb155;
e_buf = 16'h0000;
n_buf = 16'hd93c;
r_buf = 16'h26c3;
t_buf = 16'h49d7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'had4a;
e_buf = 16'h0000;
n_buf = 16'hb410;
r_buf = 16'h4bef;
t_buf = 16'h52c9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd1c2;
e_buf = 16'h0000;
n_buf = 16'h4aa2;
r_buf = 16'hb55d;
t_buf = 16'h4bc3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h33a1;
e_buf = 16'h0000;
n_buf = 16'hd92a;
r_buf = 16'h26d5;
t_buf = 16'hd4b9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he799;
e_buf = 16'h0000;
n_buf = 16'h30bb;
r_buf = 16'hcf44;
t_buf = 16'h7742;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1e70;
e_buf = 16'h0000;
n_buf = 16'hfbb2;
r_buf = 16'h044d;
t_buf = 16'h6f7d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1fed;
e_buf = 16'h0000;
n_buf = 16'h3c25;
r_buf = 16'hc3da;
t_buf = 16'ha9a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7f41;
e_buf = 16'h0000;
n_buf = 16'h9d64;
r_buf = 16'h629b;
t_buf = 16'h5e12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4993;
e_buf = 16'h0000;
n_buf = 16'he38d;
r_buf = 16'h1c72;
t_buf = 16'h4afe;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h65e0;
e_buf = 16'h0000;
n_buf = 16'h97da;
r_buf = 16'h6825;
t_buf = 16'he98f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha6e1;
e_buf = 16'h0000;
n_buf = 16'h560d;
r_buf = 16'ha9f2;
t_buf = 16'hdc90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h41a8;
e_buf = 16'h0000;
n_buf = 16'h9403;
r_buf = 16'h6bfc;
t_buf = 16'hdc64;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h278d;
e_buf = 16'h0000;
n_buf = 16'hf2e3;
r_buf = 16'h0d1c;
t_buf = 16'h2d64;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h350d;
e_buf = 16'h0000;
n_buf = 16'h64c2;
r_buf = 16'h9b3d;
t_buf = 16'h4af9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h65bf;
e_buf = 16'h0000;
n_buf = 16'h06d8;
r_buf = 16'hf927;
t_buf = 16'hc7ae;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha418;
e_buf = 16'h0000;
n_buf = 16'ha5ac;
r_buf = 16'h5a53;
t_buf = 16'h2b94;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h28b4;
e_buf = 16'h0000;
n_buf = 16'h014e;
r_buf = 16'hfeb1;
t_buf = 16'h1e9f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0ac7;
e_buf = 16'h0000;
n_buf = 16'h2b9c;
r_buf = 16'hd463;
t_buf = 16'hdd74;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0ba1;
e_buf = 16'h0000;
n_buf = 16'hfef0;
r_buf = 16'h010f;
t_buf = 16'h090e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hff3e;
e_buf = 16'h0000;
n_buf = 16'h2b28;
r_buf = 16'hd4d7;
t_buf = 16'h17df;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h985f;
e_buf = 16'h0000;
n_buf = 16'hb4d4;
r_buf = 16'h4b2b;
t_buf = 16'ha5f8;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf2ad;
e_buf = 16'h0000;
n_buf = 16'h8092;
r_buf = 16'h7f6d;
t_buf = 16'h7843;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9558;
e_buf = 16'h0000;
n_buf = 16'h90c7;
r_buf = 16'h6f38;
t_buf = 16'hc0a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcc24;
e_buf = 16'h0000;
n_buf = 16'h3a18;
r_buf = 16'hc5e7;
t_buf = 16'hcb06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hda64;
e_buf = 16'h0000;
n_buf = 16'h5ffb;
r_buf = 16'ha004;
t_buf = 16'hcfb6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3744;
e_buf = 16'h0000;
n_buf = 16'hfb69;
r_buf = 16'h0496;
t_buf = 16'h5f80;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2188;
e_buf = 16'h0000;
n_buf = 16'h324d;
r_buf = 16'hcdb2;
t_buf = 16'h1599;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9f98;
e_buf = 16'h0000;
n_buf = 16'h0326;
r_buf = 16'hfcd9;
t_buf = 16'he4e4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7cf0;
e_buf = 16'h0000;
n_buf = 16'h013d;
r_buf = 16'hfec2;
t_buf = 16'h1237;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2577;
e_buf = 16'h0000;
n_buf = 16'hc541;
r_buf = 16'h3abe;
t_buf = 16'h89fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h02ee;
e_buf = 16'h0000;
n_buf = 16'h8131;
r_buf = 16'h7ece;
t_buf = 16'h4b0f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1ac9;
e_buf = 16'h0000;
n_buf = 16'h3313;
r_buf = 16'hccec;
t_buf = 16'ha0a3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2a20;
e_buf = 16'h0000;
n_buf = 16'h5e6b;
r_buf = 16'ha194;
t_buf = 16'h9bc4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h32ae;
e_buf = 16'h0000;
n_buf = 16'h8a24;
r_buf = 16'h75db;
t_buf = 16'h1fca;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3ac1;
e_buf = 16'h0000;
n_buf = 16'hc8ce;
r_buf = 16'h3731;
t_buf = 16'hf6b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h755a;
e_buf = 16'h0000;
n_buf = 16'heb8a;
r_buf = 16'h1475;
t_buf = 16'hfb05;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3ed;
e_buf = 16'h0000;
n_buf = 16'hf364;
r_buf = 16'h0c9b;
t_buf = 16'ha19e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h60c6;
e_buf = 16'h0000;
n_buf = 16'hdc3b;
r_buf = 16'h23c4;
t_buf = 16'hc010;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9381;
e_buf = 16'h0000;
n_buf = 16'he8f8;
r_buf = 16'h1707;
t_buf = 16'h4f5f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5c94;
e_buf = 16'h0000;
n_buf = 16'h8c5f;
r_buf = 16'h73a0;
t_buf = 16'hae26;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4c3e;
e_buf = 16'h0000;
n_buf = 16'he507;
r_buf = 16'h1af8;
t_buf = 16'he824;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8be0;
e_buf = 16'h0000;
n_buf = 16'h3b6f;
r_buf = 16'hc490;
t_buf = 16'hc012;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h64b0;
e_buf = 16'h0000;
n_buf = 16'h5aa3;
r_buf = 16'ha55c;
t_buf = 16'hed41;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd3b5;
e_buf = 16'h0000;
n_buf = 16'h678a;
r_buf = 16'h9875;
t_buf = 16'hd1ae;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd974;
e_buf = 16'h0000;
n_buf = 16'h8a29;
r_buf = 16'h75d6;
t_buf = 16'h3272;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h26bd;
e_buf = 16'h0000;
n_buf = 16'h8386;
r_buf = 16'h7c79;
t_buf = 16'hc618;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha6f2;
e_buf = 16'h0000;
n_buf = 16'hf922;
r_buf = 16'h06dd;
t_buf = 16'h3810;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1ad0;
e_buf = 16'h0000;
n_buf = 16'h5804;
r_buf = 16'ha7fb;
t_buf = 16'hf2bb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc7ce;
e_buf = 16'h0000;
n_buf = 16'he711;
r_buf = 16'h18ee;
t_buf = 16'hc2b0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfd1a;
e_buf = 16'h0000;
n_buf = 16'hf3d4;
r_buf = 16'h0c2b;
t_buf = 16'hbebb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3736;
e_buf = 16'h0000;
n_buf = 16'h3418;
r_buf = 16'hcbe7;
t_buf = 16'haee5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h98a3;
e_buf = 16'h0000;
n_buf = 16'hd8f3;
r_buf = 16'h270c;
t_buf = 16'hd8e7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2e59;
e_buf = 16'h0000;
n_buf = 16'h5c4e;
r_buf = 16'ha3b1;
t_buf = 16'h0ab5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfba5;
e_buf = 16'h0000;
n_buf = 16'h93ea;
r_buf = 16'h6c15;
t_buf = 16'h4184;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1b48;
e_buf = 16'h0000;
n_buf = 16'h2cfa;
r_buf = 16'hd305;
t_buf = 16'he86e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7ce7;
e_buf = 16'h0000;
n_buf = 16'h5a70;
r_buf = 16'ha58f;
t_buf = 16'h3bf4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hacbe;
e_buf = 16'h0000;
n_buf = 16'ha82b;
r_buf = 16'h57d4;
t_buf = 16'hf521;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h25fd;
e_buf = 16'h0000;
n_buf = 16'h7589;
r_buf = 16'h8a76;
t_buf = 16'h2a57;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h053b;
e_buf = 16'h0000;
n_buf = 16'hb461;
r_buf = 16'h4b9e;
t_buf = 16'h3058;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h905c;
e_buf = 16'h0000;
n_buf = 16'he8e5;
r_buf = 16'h171a;
t_buf = 16'h79c7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8363;
e_buf = 16'h0000;
n_buf = 16'h7feb;
r_buf = 16'h8014;
t_buf = 16'ha7d5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h67e9;
e_buf = 16'h0000;
n_buf = 16'h44ef;
r_buf = 16'hbb10;
t_buf = 16'ha14e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcb01;
e_buf = 16'h0000;
n_buf = 16'h4d42;
r_buf = 16'hb2bd;
t_buf = 16'hacda;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha36b;
e_buf = 16'h0000;
n_buf = 16'ha8c2;
r_buf = 16'h573d;
t_buf = 16'h71a5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdbc8;
e_buf = 16'h0000;
n_buf = 16'h7c68;
r_buf = 16'h8397;
t_buf = 16'h7b2a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hae0f;
e_buf = 16'h0000;
n_buf = 16'h8c49;
r_buf = 16'h73b6;
t_buf = 16'ha89b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6216;
e_buf = 16'h0000;
n_buf = 16'hcecb;
r_buf = 16'h3134;
t_buf = 16'h6688;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6c59;
e_buf = 16'h0000;
n_buf = 16'h9be3;
r_buf = 16'h641c;
t_buf = 16'he227;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1a1b;
e_buf = 16'h0000;
n_buf = 16'h9285;
r_buf = 16'h6d7a;
t_buf = 16'h7c5e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he0ae;
e_buf = 16'h0000;
n_buf = 16'hf505;
r_buf = 16'h0afa;
t_buf = 16'h8dac;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3d95;
e_buf = 16'h0000;
n_buf = 16'hf87f;
r_buf = 16'h0780;
t_buf = 16'hd46c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h856f;
e_buf = 16'h0000;
n_buf = 16'hbab9;
r_buf = 16'h4546;
t_buf = 16'h4e1f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec2f;
e_buf = 16'h0000;
n_buf = 16'h2741;
r_buf = 16'hd8be;
t_buf = 16'h0035;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7ed2;
e_buf = 16'h0000;
n_buf = 16'h0176;
r_buf = 16'hfe89;
t_buf = 16'he6b1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcef3;
e_buf = 16'h0000;
n_buf = 16'h7bc7;
r_buf = 16'h8438;
t_buf = 16'hff93;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hade7;
e_buf = 16'h0000;
n_buf = 16'h6239;
r_buf = 16'h9dc6;
t_buf = 16'h7acd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9204;
e_buf = 16'h0000;
n_buf = 16'ha11b;
r_buf = 16'h5ee4;
t_buf = 16'h95c7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'heac3;
e_buf = 16'h0000;
n_buf = 16'hc89d;
r_buf = 16'h3762;
t_buf = 16'hb7d5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hac72;
e_buf = 16'h0000;
n_buf = 16'h0487;
r_buf = 16'hfb78;
t_buf = 16'h5d6a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he345;
e_buf = 16'h0000;
n_buf = 16'hdb61;
r_buf = 16'h249e;
t_buf = 16'h3560;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc241;
e_buf = 16'h0000;
n_buf = 16'h5d59;
r_buf = 16'ha2a6;
t_buf = 16'h36fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h528c;
e_buf = 16'h0000;
n_buf = 16'hd20b;
r_buf = 16'h2df4;
t_buf = 16'h1c58;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7386;
e_buf = 16'h0000;
n_buf = 16'hb337;
r_buf = 16'h4cc8;
t_buf = 16'h3895;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd562;
e_buf = 16'h0000;
n_buf = 16'hf463;
r_buf = 16'h0b9c;
t_buf = 16'h11a7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd273;
e_buf = 16'h0000;
n_buf = 16'haa37;
r_buf = 16'h55c8;
t_buf = 16'ha607;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7f99;
e_buf = 16'h0000;
n_buf = 16'he2dc;
r_buf = 16'h1d23;
t_buf = 16'h499f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec82;
e_buf = 16'h0000;
n_buf = 16'hdca7;
r_buf = 16'h2358;
t_buf = 16'hb515;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hff88;
e_buf = 16'h0000;
n_buf = 16'hf03e;
r_buf = 16'h0fc1;
t_buf = 16'h06cd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4d8a;
e_buf = 16'h0000;
n_buf = 16'ha1b7;
r_buf = 16'h5e48;
t_buf = 16'ha45d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7fa7;
e_buf = 16'h0000;
n_buf = 16'hbd91;
r_buf = 16'h426e;
t_buf = 16'h77ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9b3b;
e_buf = 16'h0000;
n_buf = 16'h3218;
r_buf = 16'hcde7;
t_buf = 16'hfdfb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha293;
e_buf = 16'h0000;
n_buf = 16'h8333;
r_buf = 16'h7ccc;
t_buf = 16'hae06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9605;
e_buf = 16'h0000;
n_buf = 16'hcae8;
r_buf = 16'h3517;
t_buf = 16'h5d01;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hab89;
e_buf = 16'h0000;
n_buf = 16'hcf23;
r_buf = 16'h30dc;
t_buf = 16'h3b71;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4623;
e_buf = 16'h0000;
n_buf = 16'h7d8f;
r_buf = 16'h8270;
t_buf = 16'h9183;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfec;
e_buf = 16'h0000;
n_buf = 16'h2116;
r_buf = 16'hdee9;
t_buf = 16'hc798;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3ce;
e_buf = 16'h0000;
n_buf = 16'h1999;
r_buf = 16'he666;
t_buf = 16'ha351;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h33b5;
e_buf = 16'h0000;
n_buf = 16'h84c8;
r_buf = 16'h7b37;
t_buf = 16'h4374;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8903;
e_buf = 16'h0000;
n_buf = 16'h8069;
r_buf = 16'h7f96;
t_buf = 16'h2722;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8af5;
e_buf = 16'h0000;
n_buf = 16'hc703;
r_buf = 16'h38fc;
t_buf = 16'hfc92;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hed34;
e_buf = 16'h0000;
n_buf = 16'h262c;
r_buf = 16'hd9d3;
t_buf = 16'hc88a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9c19;
e_buf = 16'h0000;
n_buf = 16'h8fb5;
r_buf = 16'h704a;
t_buf = 16'h22ee;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8e2f;
e_buf = 16'h0000;
n_buf = 16'hae90;
r_buf = 16'h516f;
t_buf = 16'h3683;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hee6a;
e_buf = 16'h0000;
n_buf = 16'h349a;
r_buf = 16'hcb65;
t_buf = 16'hd7c2;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8399;
e_buf = 16'h0000;
n_buf = 16'h475b;
r_buf = 16'hb8a4;
t_buf = 16'h88ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3801;
e_buf = 16'h0000;
n_buf = 16'h6d14;
r_buf = 16'h92eb;
t_buf = 16'h3d39;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h013f;
e_buf = 16'h0000;
n_buf = 16'hcd57;
r_buf = 16'h32a8;
t_buf = 16'h0175;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h027c;
e_buf = 16'h0000;
n_buf = 16'hf320;
r_buf = 16'h0cdf;
t_buf = 16'he286;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hada2;
e_buf = 16'h0000;
n_buf = 16'h18ba;
r_buf = 16'he745;
t_buf = 16'h6cfc;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5718;
e_buf = 16'h0000;
n_buf = 16'h0e5e;
r_buf = 16'hf1a1;
t_buf = 16'h20e9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hca79;
e_buf = 16'h0000;
n_buf = 16'h7d0b;
r_buf = 16'h82f4;
t_buf = 16'hdb99;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb4a1;
e_buf = 16'h0000;
n_buf = 16'h7b29;
r_buf = 16'h84d6;
t_buf = 16'h6f39;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc168;
e_buf = 16'h0000;
n_buf = 16'hfc4c;
r_buf = 16'h03b3;
t_buf = 16'hd4b7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf66a;
e_buf = 16'h0000;
n_buf = 16'hdeb8;
r_buf = 16'h2147;
t_buf = 16'h6f1c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf0bb;
e_buf = 16'h0000;
n_buf = 16'h576c;
r_buf = 16'ha893;
t_buf = 16'h9a41;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbf3d;
e_buf = 16'h0000;
n_buf = 16'h5d5f;
r_buf = 16'ha2a0;
t_buf = 16'h6732;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6403;
e_buf = 16'h0000;
n_buf = 16'h79fa;
r_buf = 16'h8605;
t_buf = 16'h8dd1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he625;
e_buf = 16'h0000;
n_buf = 16'h91eb;
r_buf = 16'h6e14;
t_buf = 16'ha366;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7350;
e_buf = 16'h0000;
n_buf = 16'h3c96;
r_buf = 16'hc369;
t_buf = 16'h8610;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5179;
e_buf = 16'h0000;
n_buf = 16'h8ded;
r_buf = 16'h7212;
t_buf = 16'hbc76;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h34ce;
e_buf = 16'h0000;
n_buf = 16'had08;
r_buf = 16'h52f7;
t_buf = 16'h2777;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd170;
e_buf = 16'h0000;
n_buf = 16'h3328;
r_buf = 16'hccd7;
t_buf = 16'h37b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1db9;
e_buf = 16'h0000;
n_buf = 16'h42f4;
r_buf = 16'hbd0b;
t_buf = 16'hdb12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5263;
e_buf = 16'h0000;
n_buf = 16'hf0e6;
r_buf = 16'h0f19;
t_buf = 16'h9409;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h72ad;
e_buf = 16'h0000;
n_buf = 16'h5c53;
r_buf = 16'ha3ac;
t_buf = 16'h7603;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0914;
e_buf = 16'h0000;
n_buf = 16'h8135;
r_buf = 16'h7eca;
t_buf = 16'hc874;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7002;
e_buf = 16'h0000;
n_buf = 16'h95dd;
r_buf = 16'h6a22;
t_buf = 16'h3bcb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h866d;
e_buf = 16'h0000;
n_buf = 16'h69d4;
r_buf = 16'h962b;
t_buf = 16'h565a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5f3d;
e_buf = 16'h0000;
n_buf = 16'h0d49;
r_buf = 16'hf2b6;
t_buf = 16'hb8f0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h25fb;
e_buf = 16'h0000;
n_buf = 16'h7c24;
r_buf = 16'h83db;
t_buf = 16'h9544;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2281;
e_buf = 16'h0000;
n_buf = 16'hcdff;
r_buf = 16'h3200;
t_buf = 16'hc2b6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfde;
e_buf = 16'h0000;
n_buf = 16'hd037;
r_buf = 16'h2fc8;
t_buf = 16'h713b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0359;
e_buf = 16'h0000;
n_buf = 16'h9643;
r_buf = 16'h69bc;
t_buf = 16'h99d4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h41c3;
e_buf = 16'h0000;
n_buf = 16'h5b56;
r_buf = 16'ha4a9;
t_buf = 16'h11f4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1f7a;
e_buf = 16'h0000;
n_buf = 16'hb9af;
r_buf = 16'h4650;
t_buf = 16'hefe9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9a43;
e_buf = 16'h0000;
n_buf = 16'h6a17;
r_buf = 16'h95e8;
t_buf = 16'hfb94;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h23fb;
e_buf = 16'h0000;
n_buf = 16'h9008;
r_buf = 16'h6ff7;
t_buf = 16'hc724;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc8bf;
e_buf = 16'h0000;
n_buf = 16'h5898;
r_buf = 16'ha767;
t_buf = 16'hfc15;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h69e2;
e_buf = 16'h0000;
n_buf = 16'hdba8;
r_buf = 16'h2457;
t_buf = 16'h088f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h27e9;
e_buf = 16'h0000;
n_buf = 16'h0067;
r_buf = 16'hff98;
t_buf = 16'h3c4a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h283c;
e_buf = 16'h0000;
n_buf = 16'hbf02;
r_buf = 16'h40fd;
t_buf = 16'haa15;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd7a3;
e_buf = 16'h0000;
n_buf = 16'h89d9;
r_buf = 16'h7626;
t_buf = 16'hb031;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7a8c;
e_buf = 16'h0000;
n_buf = 16'h9ebe;
r_buf = 16'h6141;
t_buf = 16'ha21e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6106;
e_buf = 16'h0000;
n_buf = 16'h8a44;
r_buf = 16'h75bb;
t_buf = 16'hebaf;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h178e;
e_buf = 16'h0000;
n_buf = 16'h0129;
r_buf = 16'hfed6;
t_buf = 16'h5b17;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h953c;
e_buf = 16'h0000;
n_buf = 16'h9f9d;
r_buf = 16'h6062;
t_buf = 16'h26e9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha436;
e_buf = 16'h0000;
n_buf = 16'h6b43;
r_buf = 16'h94bc;
t_buf = 16'h46c0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4b5c;
e_buf = 16'h0000;
n_buf = 16'hc954;
r_buf = 16'h36ab;
t_buf = 16'h578e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h79cc;
e_buf = 16'h0000;
n_buf = 16'haf4e;
r_buf = 16'h50b1;
t_buf = 16'h9120;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb7d7;
e_buf = 16'h0000;
n_buf = 16'h9cc9;
r_buf = 16'h6336;
t_buf = 16'h94fb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfcc;
e_buf = 16'h0000;
n_buf = 16'h6c9a;
r_buf = 16'h9365;
t_buf = 16'h516a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb4d4;
e_buf = 16'h0000;
n_buf = 16'h54c5;
r_buf = 16'hab3a;
t_buf = 16'hc95f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2e70;
e_buf = 16'h0000;
n_buf = 16'h1bc3;
r_buf = 16'he43c;
t_buf = 16'ha743;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hce9b;
e_buf = 16'h0000;
n_buf = 16'h7549;
r_buf = 16'h8ab6;
t_buf = 16'h5a43;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h30ef;
e_buf = 16'h0000;
n_buf = 16'h1c04;
r_buf = 16'he3fb;
t_buf = 16'h9a28;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h786e;
e_buf = 16'h0000;
n_buf = 16'h9990;
r_buf = 16'h666f;
t_buf = 16'h3a9a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he97d;
e_buf = 16'h0000;
n_buf = 16'h5e42;
r_buf = 16'ha1bd;
t_buf = 16'h3152;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h10fc;
e_buf = 16'h0000;
n_buf = 16'h0729;
r_buf = 16'hf8d6;
t_buf = 16'h4a11;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3ff7;
e_buf = 16'h0000;
n_buf = 16'h4404;
r_buf = 16'hbbfb;
t_buf = 16'h626f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hccc9;
e_buf = 16'h0000;
n_buf = 16'hcdf8;
r_buf = 16'h3207;
t_buf = 16'h958f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2c21;
e_buf = 16'h0000;
n_buf = 16'h652c;
r_buf = 16'h9ad3;
t_buf = 16'hbbc4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h15ab;
e_buf = 16'h0000;
n_buf = 16'h3ac7;
r_buf = 16'hc538;
t_buf = 16'hd03f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2a7d;
e_buf = 16'h0000;
n_buf = 16'hae1f;
r_buf = 16'h51e0;
t_buf = 16'ha87c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h843b;
e_buf = 16'h0000;
n_buf = 16'ha2a7;
r_buf = 16'h5d58;
t_buf = 16'h7d90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec4b;
e_buf = 16'h0000;
n_buf = 16'hb79b;
r_buf = 16'h4864;
t_buf = 16'hb1b9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hde6f;
e_buf = 16'h0000;
n_buf = 16'h2d5d;
r_buf = 16'hd2a2;
t_buf = 16'ha48b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h24b6;
e_buf = 16'h0000;
n_buf = 16'h5cd1;
r_buf = 16'ha32e;
t_buf = 16'he73a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hea5f;
e_buf = 16'h0000;
n_buf = 16'h8cfe;
r_buf = 16'h7301;
t_buf = 16'hde0a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h27f7;
e_buf = 16'h0000;
n_buf = 16'h3a51;
r_buf = 16'hc5ae;
t_buf = 16'h68a6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0a17;
e_buf = 16'h0000;
n_buf = 16'h959f;
r_buf = 16'h6a60;
t_buf = 16'h191b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9eee;
e_buf = 16'h0000;
n_buf = 16'hdc0e;
r_buf = 16'h23f1;
t_buf = 16'h6229;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h10fc;
e_buf = 16'h0000;
n_buf = 16'h2e47;
r_buf = 16'hd1b8;
t_buf = 16'h1b9e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8a8f;
e_buf = 16'h0000;
n_buf = 16'h13ab;
r_buf = 16'hec54;
t_buf = 16'h1b92;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h399f;
e_buf = 16'h0000;
n_buf = 16'hdc6b;
r_buf = 16'h2394;
t_buf = 16'h1c90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1081;
e_buf = 16'h0000;
n_buf = 16'h308c;
r_buf = 16'hcf73;
t_buf = 16'h28b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2168;
e_buf = 16'h0000;
n_buf = 16'h1773;
r_buf = 16'he88c;
t_buf = 16'h17f3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdc4e;
e_buf = 16'h0000;
n_buf = 16'h7e97;
r_buf = 16'h8168;
t_buf = 16'hfa69;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0a66;
e_buf = 16'h0000;
n_buf = 16'hcc66;
r_buf = 16'h3399;
t_buf = 16'hc788;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2df0;
e_buf = 16'h0000;
n_buf = 16'h3ed3;
r_buf = 16'hc12c;
t_buf = 16'hcd53;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4cea;
e_buf = 16'h0000;
n_buf = 16'h8d10;
r_buf = 16'h72ef;
t_buf = 16'h6482;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hba02;
e_buf = 16'h0000;
n_buf = 16'h95ee;
r_buf = 16'h6a11;
t_buf = 16'hcd0d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h03e9;
e_buf = 16'h0000;
n_buf = 16'hcc0e;
r_buf = 16'h33f1;
t_buf = 16'h84ee;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2fd6;
e_buf = 16'h0000;
n_buf = 16'h17e3;
r_buf = 16'he81c;
t_buf = 16'ha5e6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc247;
e_buf = 16'h0000;
n_buf = 16'hd9ed;
r_buf = 16'h2612;
t_buf = 16'h1b98;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6a1c;
e_buf = 16'h0000;
n_buf = 16'h0a15;
r_buf = 16'hf5ea;
t_buf = 16'h588c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd80d;
e_buf = 16'h0000;
n_buf = 16'hd102;
r_buf = 16'h2efd;
t_buf = 16'hd58c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbc20;
e_buf = 16'h0000;
n_buf = 16'hbdb6;
r_buf = 16'h4249;
t_buf = 16'hcb70;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h72d6;
e_buf = 16'h0000;
n_buf = 16'hee52;
r_buf = 16'h11ad;
t_buf = 16'h6748;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd505;
e_buf = 16'h0000;
n_buf = 16'hf341;
r_buf = 16'h0cbe;
t_buf = 16'h394a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h54a1;
e_buf = 16'h0000;
n_buf = 16'h415a;
r_buf = 16'hbea5;
t_buf = 16'h2a7c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb353;
e_buf = 16'h0000;
n_buf = 16'h3dd6;
r_buf = 16'hc229;
t_buf = 16'hae09;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdca5;
e_buf = 16'h0000;
n_buf = 16'h084f;
r_buf = 16'hf7b0;
t_buf = 16'h9518;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfbd8;
e_buf = 16'h0000;
n_buf = 16'h96c0;
r_buf = 16'h693f;
t_buf = 16'hb8ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2922;
e_buf = 16'h0000;
n_buf = 16'hd77c;
r_buf = 16'h2883;
t_buf = 16'h0a12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h19ab;
e_buf = 16'h0000;
n_buf = 16'hd1ee;
r_buf = 16'h2e11;
t_buf = 16'hb144;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hccf7;
e_buf = 16'h0000;
n_buf = 16'hf18d;
r_buf = 16'h0e72;
t_buf = 16'h3ef4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h08b9;
e_buf = 16'h0000;
n_buf = 16'h2b01;
r_buf = 16'hd4fe;
t_buf = 16'h5da4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2619;
e_buf = 16'h0000;
n_buf = 16'hac51;
r_buf = 16'h53ae;
t_buf = 16'h3ca9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd43f;
e_buf = 16'h0000;
n_buf = 16'h3d26;
r_buf = 16'hc2d9;
t_buf = 16'h37fa;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hde62;
e_buf = 16'h0000;
n_buf = 16'h1209;
r_buf = 16'hedf6;
t_buf = 16'h6e66;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h195c;
e_buf = 16'h0000;
n_buf = 16'hd512;
r_buf = 16'h2aed;
t_buf = 16'h64a8;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha7f5;
e_buf = 16'h0000;
n_buf = 16'h154e;
r_buf = 16'heab1;
t_buf = 16'h22a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbc20;
e_buf = 16'h0000;
n_buf = 16'h5db5;
r_buf = 16'ha24a;
t_buf = 16'h9179;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h75f2;
e_buf = 16'h0000;
n_buf = 16'hde3a;
r_buf = 16'h21c5;
t_buf = 16'h07c9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0e7f;
e_buf = 16'h0000;
n_buf = 16'hd656;
r_buf = 16'h29a9;
t_buf = 16'h295f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf7f6;
e_buf = 16'h0000;
n_buf = 16'h0445;
r_buf = 16'hfbba;
t_buf = 16'hf135;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf320;
e_buf = 16'h0000;
n_buf = 16'hba8e;
r_buf = 16'h4571;
t_buf = 16'h6470;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5f0e;
e_buf = 16'h0000;
n_buf = 16'h73f7;
r_buf = 16'h8c08;
t_buf = 16'hf206;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha8f4;
e_buf = 16'h0000;
n_buf = 16'h33db;
r_buf = 16'hcc24;
t_buf = 16'ha4fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8147;
e_buf = 16'h0000;
n_buf = 16'h03ba;
r_buf = 16'hfc45;
t_buf = 16'hd8ed;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfe39;
e_buf = 16'h0000;
n_buf = 16'haa40;
r_buf = 16'h55bf;
t_buf = 16'h062b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h61d9;
e_buf = 16'h0000;
n_buf = 16'hc10f;
r_buf = 16'h3ef0;
t_buf = 16'h9d89;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdd9e;
e_buf = 16'h0000;
n_buf = 16'h2284;
r_buf = 16'hdd7b;
t_buf = 16'h8f40;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he6ad;
e_buf = 16'h0000;
n_buf = 16'hc16e;
r_buf = 16'h3e91;
t_buf = 16'hd5f5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h798f;
e_buf = 16'h0000;
n_buf = 16'h816a;
r_buf = 16'h7e95;
t_buf = 16'h23da;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h87a1;
e_buf = 16'h0000;
n_buf = 16'h47fc;
r_buf = 16'hb803;
t_buf = 16'h7185;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2923;
e_buf = 16'h0000;
n_buf = 16'h1d03;
r_buf = 16'he2fc;
t_buf = 16'hfa46;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h809f;
e_buf = 16'h0000;
n_buf = 16'h3fe3;
r_buf = 16'hc01c;
t_buf = 16'had98;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9850;
e_buf = 16'h0000;
n_buf = 16'hb476;
r_buf = 16'h4b89;
t_buf = 16'h1965;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h044d;
e_buf = 16'h0000;
n_buf = 16'h84c5;
r_buf = 16'h7b3a;
t_buf = 16'h149c;
nprime0_buf = 16'h0000;


	#3000
	startCompute = 1;
	#10
	startCompute = 0;


#10000000
getResult = 1;
#10
getResult = 0;

#1000
reset = 1;
startInput = 0;
#10
reset = 0;
#100 
startInput = 1;	


#10
m_buf = 16'h6d1d;
e_buf = 16'h000f;
n_buf = 16'h898f;
r_buf = 16'h7671;
t_buf = 16'h289e;
nprime0_buf = 16'h8a91;
#10
m_buf = 16'h42cb;
e_buf = 16'h0000;
n_buf = 16'h5fec;
r_buf = 16'ha013;
t_buf = 16'hacaa;
nprime0_buf = 16'ha3b1;
#10
m_buf = 16'h8051;
e_buf = 16'h0000;
n_buf = 16'hbd79;
r_buf = 16'h4286;
t_buf = 16'h3f82;
nprime0_buf = 16'h2df6;
#10
m_buf = 16'h95d1;
e_buf = 16'h0000;
n_buf = 16'h1622;
r_buf = 16'he9dd;
t_buf = 16'h7305;
nprime0_buf = 16'h3bea;
#10
m_buf = 16'h0933;
e_buf = 16'h0000;
n_buf = 16'hca16;
r_buf = 16'h35e9;
t_buf = 16'hf2c5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc6f0;
e_buf = 16'h0000;
n_buf = 16'h705f;
r_buf = 16'h8fa0;
t_buf = 16'h2b90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0f4e;
e_buf = 16'h0000;
n_buf = 16'h0806;
r_buf = 16'hf7f9;
t_buf = 16'h6657;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2aa5;
e_buf = 16'h0000;
n_buf = 16'ha9ec;
r_buf = 16'h5613;
t_buf = 16'h4906;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8043;
e_buf = 16'h0000;
n_buf = 16'h3d15;
r_buf = 16'hc2ea;
t_buf = 16'h0a06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6e64;
e_buf = 16'h0000;
n_buf = 16'h8228;
r_buf = 16'h7dd7;
t_buf = 16'h0040;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4efe;
e_buf = 16'h0000;
n_buf = 16'h6215;
r_buf = 16'h9dea;
t_buf = 16'h0115;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3123;
e_buf = 16'h0000;
n_buf = 16'h1ba1;
r_buf = 16'he45e;
t_buf = 16'h41d7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfdeb;
e_buf = 16'h0000;
n_buf = 16'h03e3;
r_buf = 16'hfc1c;
t_buf = 16'h4bdb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5bc7;
e_buf = 16'h0000;
n_buf = 16'hc748;
r_buf = 16'h38b7;
t_buf = 16'hd1a3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h73e5;
e_buf = 16'h0000;
n_buf = 16'h21a4;
r_buf = 16'hde5b;
t_buf = 16'hb841;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1d71;
e_buf = 16'h0000;
n_buf = 16'h29e8;
r_buf = 16'hd617;
t_buf = 16'h4255;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfe8c;
e_buf = 16'h0000;
n_buf = 16'h3844;
r_buf = 16'hc7bb;
t_buf = 16'h73e0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1058;
e_buf = 16'h0000;
n_buf = 16'h855c;
r_buf = 16'h7aa3;
t_buf = 16'hdf44;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5396;
e_buf = 16'h0000;
n_buf = 16'h107e;
r_buf = 16'hef81;
t_buf = 16'hbcdf;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd26d;
e_buf = 16'h0000;
n_buf = 16'hd707;
r_buf = 16'h28f8;
t_buf = 16'h0d21;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8266;
e_buf = 16'h0000;
n_buf = 16'h5db9;
r_buf = 16'ha246;
t_buf = 16'hfa55;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdd13;
e_buf = 16'h0000;
n_buf = 16'h64ac;
r_buf = 16'h9b53;
t_buf = 16'h386e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf267;
e_buf = 16'h0000;
n_buf = 16'h92d8;
r_buf = 16'h6d27;
t_buf = 16'hce5f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hda54;
e_buf = 16'h0000;
n_buf = 16'h5eda;
r_buf = 16'ha125;
t_buf = 16'hef79;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8b57;
e_buf = 16'h0000;
n_buf = 16'h8dfc;
r_buf = 16'h7203;
t_buf = 16'h8c2e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3b6;
e_buf = 16'h0000;
n_buf = 16'h7d5c;
r_buf = 16'h82a3;
t_buf = 16'h2b88;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0911;
e_buf = 16'h0000;
n_buf = 16'h8a43;
r_buf = 16'h75bc;
t_buf = 16'hbaa2;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0712;
e_buf = 16'h0000;
n_buf = 16'hbb96;
r_buf = 16'h4469;
t_buf = 16'ha401;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb5b7;
e_buf = 16'h0000;
n_buf = 16'h3986;
r_buf = 16'hc679;
t_buf = 16'hf001;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he72b;
e_buf = 16'h0000;
n_buf = 16'h0792;
r_buf = 16'hf86d;
t_buf = 16'h0135;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdbd2;
e_buf = 16'h0000;
n_buf = 16'h5d68;
r_buf = 16'ha297;
t_buf = 16'h1e91;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h869b;
e_buf = 16'h0000;
n_buf = 16'h7825;
r_buf = 16'h87da;
t_buf = 16'h432c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd488;
e_buf = 16'h0000;
n_buf = 16'hfbac;
r_buf = 16'h0453;
t_buf = 16'hd484;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h739c;
e_buf = 16'h0000;
n_buf = 16'h0b21;
r_buf = 16'hf4de;
t_buf = 16'h9f25;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcd8f;
e_buf = 16'h0000;
n_buf = 16'hc8d6;
r_buf = 16'h3729;
t_buf = 16'h6bf1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc09f;
e_buf = 16'h0000;
n_buf = 16'h4efb;
r_buf = 16'hb104;
t_buf = 16'h192d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb155;
e_buf = 16'h0000;
n_buf = 16'hd93c;
r_buf = 16'h26c3;
t_buf = 16'h49d7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'had4a;
e_buf = 16'h0000;
n_buf = 16'hb410;
r_buf = 16'h4bef;
t_buf = 16'h52c9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd1c2;
e_buf = 16'h0000;
n_buf = 16'h4aa2;
r_buf = 16'hb55d;
t_buf = 16'h4bc3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h33a1;
e_buf = 16'h0000;
n_buf = 16'hd92a;
r_buf = 16'h26d5;
t_buf = 16'hd4b9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he799;
e_buf = 16'h0000;
n_buf = 16'h30bb;
r_buf = 16'hcf44;
t_buf = 16'h7742;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1e70;
e_buf = 16'h0000;
n_buf = 16'hfbb2;
r_buf = 16'h044d;
t_buf = 16'h6f7d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1fed;
e_buf = 16'h0000;
n_buf = 16'h3c25;
r_buf = 16'hc3da;
t_buf = 16'ha9a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7f41;
e_buf = 16'h0000;
n_buf = 16'h9d64;
r_buf = 16'h629b;
t_buf = 16'h5e12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4993;
e_buf = 16'h0000;
n_buf = 16'he38d;
r_buf = 16'h1c72;
t_buf = 16'h4afe;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h65e0;
e_buf = 16'h0000;
n_buf = 16'h97da;
r_buf = 16'h6825;
t_buf = 16'he98f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha6e1;
e_buf = 16'h0000;
n_buf = 16'h560d;
r_buf = 16'ha9f2;
t_buf = 16'hdc90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h41a8;
e_buf = 16'h0000;
n_buf = 16'h9403;
r_buf = 16'h6bfc;
t_buf = 16'hdc64;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h278d;
e_buf = 16'h0000;
n_buf = 16'hf2e3;
r_buf = 16'h0d1c;
t_buf = 16'h2d64;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h350d;
e_buf = 16'h0000;
n_buf = 16'h64c2;
r_buf = 16'h9b3d;
t_buf = 16'h4af9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h65bf;
e_buf = 16'h0000;
n_buf = 16'h06d8;
r_buf = 16'hf927;
t_buf = 16'hc7ae;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha418;
e_buf = 16'h0000;
n_buf = 16'ha5ac;
r_buf = 16'h5a53;
t_buf = 16'h2b94;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h28b4;
e_buf = 16'h0000;
n_buf = 16'h014e;
r_buf = 16'hfeb1;
t_buf = 16'h1e9f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0ac7;
e_buf = 16'h0000;
n_buf = 16'h2b9c;
r_buf = 16'hd463;
t_buf = 16'hdd74;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0ba1;
e_buf = 16'h0000;
n_buf = 16'hfef0;
r_buf = 16'h010f;
t_buf = 16'h090e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hff3e;
e_buf = 16'h0000;
n_buf = 16'h2b28;
r_buf = 16'hd4d7;
t_buf = 16'h17df;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h985f;
e_buf = 16'h0000;
n_buf = 16'hb4d4;
r_buf = 16'h4b2b;
t_buf = 16'ha5f8;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf2ad;
e_buf = 16'h0000;
n_buf = 16'h8092;
r_buf = 16'h7f6d;
t_buf = 16'h7843;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9558;
e_buf = 16'h0000;
n_buf = 16'h90c7;
r_buf = 16'h6f38;
t_buf = 16'hc0a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcc24;
e_buf = 16'h0000;
n_buf = 16'h3a18;
r_buf = 16'hc5e7;
t_buf = 16'hcb06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hda64;
e_buf = 16'h0000;
n_buf = 16'h5ffb;
r_buf = 16'ha004;
t_buf = 16'hcfb6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3744;
e_buf = 16'h0000;
n_buf = 16'hfb69;
r_buf = 16'h0496;
t_buf = 16'h5f80;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2188;
e_buf = 16'h0000;
n_buf = 16'h324d;
r_buf = 16'hcdb2;
t_buf = 16'h1599;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9f98;
e_buf = 16'h0000;
n_buf = 16'h0326;
r_buf = 16'hfcd9;
t_buf = 16'he4e4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7cf0;
e_buf = 16'h0000;
n_buf = 16'h013d;
r_buf = 16'hfec2;
t_buf = 16'h1237;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2577;
e_buf = 16'h0000;
n_buf = 16'hc541;
r_buf = 16'h3abe;
t_buf = 16'h89fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h02ee;
e_buf = 16'h0000;
n_buf = 16'h8131;
r_buf = 16'h7ece;
t_buf = 16'h4b0f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1ac9;
e_buf = 16'h0000;
n_buf = 16'h3313;
r_buf = 16'hccec;
t_buf = 16'ha0a3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2a20;
e_buf = 16'h0000;
n_buf = 16'h5e6b;
r_buf = 16'ha194;
t_buf = 16'h9bc4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h32ae;
e_buf = 16'h0000;
n_buf = 16'h8a24;
r_buf = 16'h75db;
t_buf = 16'h1fca;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3ac1;
e_buf = 16'h0000;
n_buf = 16'hc8ce;
r_buf = 16'h3731;
t_buf = 16'hf6b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h755a;
e_buf = 16'h0000;
n_buf = 16'heb8a;
r_buf = 16'h1475;
t_buf = 16'hfb05;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3ed;
e_buf = 16'h0000;
n_buf = 16'hf364;
r_buf = 16'h0c9b;
t_buf = 16'ha19e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h60c6;
e_buf = 16'h0000;
n_buf = 16'hdc3b;
r_buf = 16'h23c4;
t_buf = 16'hc010;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9381;
e_buf = 16'h0000;
n_buf = 16'he8f8;
r_buf = 16'h1707;
t_buf = 16'h4f5f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5c94;
e_buf = 16'h0000;
n_buf = 16'h8c5f;
r_buf = 16'h73a0;
t_buf = 16'hae26;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4c3e;
e_buf = 16'h0000;
n_buf = 16'he507;
r_buf = 16'h1af8;
t_buf = 16'he824;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8be0;
e_buf = 16'h0000;
n_buf = 16'h3b6f;
r_buf = 16'hc490;
t_buf = 16'hc012;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h64b0;
e_buf = 16'h0000;
n_buf = 16'h5aa3;
r_buf = 16'ha55c;
t_buf = 16'hed41;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd3b5;
e_buf = 16'h0000;
n_buf = 16'h678a;
r_buf = 16'h9875;
t_buf = 16'hd1ae;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd974;
e_buf = 16'h0000;
n_buf = 16'h8a29;
r_buf = 16'h75d6;
t_buf = 16'h3272;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h26bd;
e_buf = 16'h0000;
n_buf = 16'h8386;
r_buf = 16'h7c79;
t_buf = 16'hc618;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha6f2;
e_buf = 16'h0000;
n_buf = 16'hf922;
r_buf = 16'h06dd;
t_buf = 16'h3810;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1ad0;
e_buf = 16'h0000;
n_buf = 16'h5804;
r_buf = 16'ha7fb;
t_buf = 16'hf2bb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc7ce;
e_buf = 16'h0000;
n_buf = 16'he711;
r_buf = 16'h18ee;
t_buf = 16'hc2b0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfd1a;
e_buf = 16'h0000;
n_buf = 16'hf3d4;
r_buf = 16'h0c2b;
t_buf = 16'hbebb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3736;
e_buf = 16'h0000;
n_buf = 16'h3418;
r_buf = 16'hcbe7;
t_buf = 16'haee5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h98a3;
e_buf = 16'h0000;
n_buf = 16'hd8f3;
r_buf = 16'h270c;
t_buf = 16'hd8e7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2e59;
e_buf = 16'h0000;
n_buf = 16'h5c4e;
r_buf = 16'ha3b1;
t_buf = 16'h0ab5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfba5;
e_buf = 16'h0000;
n_buf = 16'h93ea;
r_buf = 16'h6c15;
t_buf = 16'h4184;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1b48;
e_buf = 16'h0000;
n_buf = 16'h2cfa;
r_buf = 16'hd305;
t_buf = 16'he86e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7ce7;
e_buf = 16'h0000;
n_buf = 16'h5a70;
r_buf = 16'ha58f;
t_buf = 16'h3bf4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hacbe;
e_buf = 16'h0000;
n_buf = 16'ha82b;
r_buf = 16'h57d4;
t_buf = 16'hf521;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h25fd;
e_buf = 16'h0000;
n_buf = 16'h7589;
r_buf = 16'h8a76;
t_buf = 16'h2a57;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h053b;
e_buf = 16'h0000;
n_buf = 16'hb461;
r_buf = 16'h4b9e;
t_buf = 16'h3058;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h905c;
e_buf = 16'h0000;
n_buf = 16'he8e5;
r_buf = 16'h171a;
t_buf = 16'h79c7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8363;
e_buf = 16'h0000;
n_buf = 16'h7feb;
r_buf = 16'h8014;
t_buf = 16'ha7d5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h67e9;
e_buf = 16'h0000;
n_buf = 16'h44ef;
r_buf = 16'hbb10;
t_buf = 16'ha14e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcb01;
e_buf = 16'h0000;
n_buf = 16'h4d42;
r_buf = 16'hb2bd;
t_buf = 16'hacda;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha36b;
e_buf = 16'h0000;
n_buf = 16'ha8c2;
r_buf = 16'h573d;
t_buf = 16'h71a5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdbc8;
e_buf = 16'h0000;
n_buf = 16'h7c68;
r_buf = 16'h8397;
t_buf = 16'h7b2a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hae0f;
e_buf = 16'h0000;
n_buf = 16'h8c49;
r_buf = 16'h73b6;
t_buf = 16'ha89b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6216;
e_buf = 16'h0000;
n_buf = 16'hcecb;
r_buf = 16'h3134;
t_buf = 16'h6688;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6c59;
e_buf = 16'h0000;
n_buf = 16'h9be3;
r_buf = 16'h641c;
t_buf = 16'he227;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1a1b;
e_buf = 16'h0000;
n_buf = 16'h9285;
r_buf = 16'h6d7a;
t_buf = 16'h7c5e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he0ae;
e_buf = 16'h0000;
n_buf = 16'hf505;
r_buf = 16'h0afa;
t_buf = 16'h8dac;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3d95;
e_buf = 16'h0000;
n_buf = 16'hf87f;
r_buf = 16'h0780;
t_buf = 16'hd46c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h856f;
e_buf = 16'h0000;
n_buf = 16'hbab9;
r_buf = 16'h4546;
t_buf = 16'h4e1f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec2f;
e_buf = 16'h0000;
n_buf = 16'h2741;
r_buf = 16'hd8be;
t_buf = 16'h0035;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7ed2;
e_buf = 16'h0000;
n_buf = 16'h0176;
r_buf = 16'hfe89;
t_buf = 16'he6b1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hcef3;
e_buf = 16'h0000;
n_buf = 16'h7bc7;
r_buf = 16'h8438;
t_buf = 16'hff93;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hade7;
e_buf = 16'h0000;
n_buf = 16'h6239;
r_buf = 16'h9dc6;
t_buf = 16'h7acd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9204;
e_buf = 16'h0000;
n_buf = 16'ha11b;
r_buf = 16'h5ee4;
t_buf = 16'h95c7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'heac3;
e_buf = 16'h0000;
n_buf = 16'hc89d;
r_buf = 16'h3762;
t_buf = 16'hb7d5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hac72;
e_buf = 16'h0000;
n_buf = 16'h0487;
r_buf = 16'hfb78;
t_buf = 16'h5d6a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he345;
e_buf = 16'h0000;
n_buf = 16'hdb61;
r_buf = 16'h249e;
t_buf = 16'h3560;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc241;
e_buf = 16'h0000;
n_buf = 16'h5d59;
r_buf = 16'ha2a6;
t_buf = 16'h36fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h528c;
e_buf = 16'h0000;
n_buf = 16'hd20b;
r_buf = 16'h2df4;
t_buf = 16'h1c58;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7386;
e_buf = 16'h0000;
n_buf = 16'hb337;
r_buf = 16'h4cc8;
t_buf = 16'h3895;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd562;
e_buf = 16'h0000;
n_buf = 16'hf463;
r_buf = 16'h0b9c;
t_buf = 16'h11a7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd273;
e_buf = 16'h0000;
n_buf = 16'haa37;
r_buf = 16'h55c8;
t_buf = 16'ha607;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7f99;
e_buf = 16'h0000;
n_buf = 16'he2dc;
r_buf = 16'h1d23;
t_buf = 16'h499f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec82;
e_buf = 16'h0000;
n_buf = 16'hdca7;
r_buf = 16'h2358;
t_buf = 16'hb515;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hff88;
e_buf = 16'h0000;
n_buf = 16'hf03e;
r_buf = 16'h0fc1;
t_buf = 16'h06cd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4d8a;
e_buf = 16'h0000;
n_buf = 16'ha1b7;
r_buf = 16'h5e48;
t_buf = 16'ha45d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7fa7;
e_buf = 16'h0000;
n_buf = 16'hbd91;
r_buf = 16'h426e;
t_buf = 16'h77ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9b3b;
e_buf = 16'h0000;
n_buf = 16'h3218;
r_buf = 16'hcde7;
t_buf = 16'hfdfb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha293;
e_buf = 16'h0000;
n_buf = 16'h8333;
r_buf = 16'h7ccc;
t_buf = 16'hae06;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9605;
e_buf = 16'h0000;
n_buf = 16'hcae8;
r_buf = 16'h3517;
t_buf = 16'h5d01;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hab89;
e_buf = 16'h0000;
n_buf = 16'hcf23;
r_buf = 16'h30dc;
t_buf = 16'h3b71;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4623;
e_buf = 16'h0000;
n_buf = 16'h7d8f;
r_buf = 16'h8270;
t_buf = 16'h9183;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfec;
e_buf = 16'h0000;
n_buf = 16'h2116;
r_buf = 16'hdee9;
t_buf = 16'hc798;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb3ce;
e_buf = 16'h0000;
n_buf = 16'h1999;
r_buf = 16'he666;
t_buf = 16'ha351;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h33b5;
e_buf = 16'h0000;
n_buf = 16'h84c8;
r_buf = 16'h7b37;
t_buf = 16'h4374;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8903;
e_buf = 16'h0000;
n_buf = 16'h8069;
r_buf = 16'h7f96;
t_buf = 16'h2722;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8af5;
e_buf = 16'h0000;
n_buf = 16'hc703;
r_buf = 16'h38fc;
t_buf = 16'hfc92;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hed34;
e_buf = 16'h0000;
n_buf = 16'h262c;
r_buf = 16'hd9d3;
t_buf = 16'hc88a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9c19;
e_buf = 16'h0000;
n_buf = 16'h8fb5;
r_buf = 16'h704a;
t_buf = 16'h22ee;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8e2f;
e_buf = 16'h0000;
n_buf = 16'hae90;
r_buf = 16'h516f;
t_buf = 16'h3683;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hee6a;
e_buf = 16'h0000;
n_buf = 16'h349a;
r_buf = 16'hcb65;
t_buf = 16'hd7c2;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8399;
e_buf = 16'h0000;
n_buf = 16'h475b;
r_buf = 16'hb8a4;
t_buf = 16'h88ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3801;
e_buf = 16'h0000;
n_buf = 16'h6d14;
r_buf = 16'h92eb;
t_buf = 16'h3d39;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h013f;
e_buf = 16'h0000;
n_buf = 16'hcd57;
r_buf = 16'h32a8;
t_buf = 16'h0175;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h027c;
e_buf = 16'h0000;
n_buf = 16'hf320;
r_buf = 16'h0cdf;
t_buf = 16'he286;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hada2;
e_buf = 16'h0000;
n_buf = 16'h18ba;
r_buf = 16'he745;
t_buf = 16'h6cfc;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5718;
e_buf = 16'h0000;
n_buf = 16'h0e5e;
r_buf = 16'hf1a1;
t_buf = 16'h20e9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hca79;
e_buf = 16'h0000;
n_buf = 16'h7d0b;
r_buf = 16'h82f4;
t_buf = 16'hdb99;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb4a1;
e_buf = 16'h0000;
n_buf = 16'h7b29;
r_buf = 16'h84d6;
t_buf = 16'h6f39;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc168;
e_buf = 16'h0000;
n_buf = 16'hfc4c;
r_buf = 16'h03b3;
t_buf = 16'hd4b7;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf66a;
e_buf = 16'h0000;
n_buf = 16'hdeb8;
r_buf = 16'h2147;
t_buf = 16'h6f1c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf0bb;
e_buf = 16'h0000;
n_buf = 16'h576c;
r_buf = 16'ha893;
t_buf = 16'h9a41;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbf3d;
e_buf = 16'h0000;
n_buf = 16'h5d5f;
r_buf = 16'ha2a0;
t_buf = 16'h6732;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6403;
e_buf = 16'h0000;
n_buf = 16'h79fa;
r_buf = 16'h8605;
t_buf = 16'h8dd1;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he625;
e_buf = 16'h0000;
n_buf = 16'h91eb;
r_buf = 16'h6e14;
t_buf = 16'ha366;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7350;
e_buf = 16'h0000;
n_buf = 16'h3c96;
r_buf = 16'hc369;
t_buf = 16'h8610;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5179;
e_buf = 16'h0000;
n_buf = 16'h8ded;
r_buf = 16'h7212;
t_buf = 16'hbc76;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h34ce;
e_buf = 16'h0000;
n_buf = 16'had08;
r_buf = 16'h52f7;
t_buf = 16'h2777;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd170;
e_buf = 16'h0000;
n_buf = 16'h3328;
r_buf = 16'hccd7;
t_buf = 16'h37b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1db9;
e_buf = 16'h0000;
n_buf = 16'h42f4;
r_buf = 16'hbd0b;
t_buf = 16'hdb12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5263;
e_buf = 16'h0000;
n_buf = 16'hf0e6;
r_buf = 16'h0f19;
t_buf = 16'h9409;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h72ad;
e_buf = 16'h0000;
n_buf = 16'h5c53;
r_buf = 16'ha3ac;
t_buf = 16'h7603;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0914;
e_buf = 16'h0000;
n_buf = 16'h8135;
r_buf = 16'h7eca;
t_buf = 16'hc874;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7002;
e_buf = 16'h0000;
n_buf = 16'h95dd;
r_buf = 16'h6a22;
t_buf = 16'h3bcb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h866d;
e_buf = 16'h0000;
n_buf = 16'h69d4;
r_buf = 16'h962b;
t_buf = 16'h565a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5f3d;
e_buf = 16'h0000;
n_buf = 16'h0d49;
r_buf = 16'hf2b6;
t_buf = 16'hb8f0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h25fb;
e_buf = 16'h0000;
n_buf = 16'h7c24;
r_buf = 16'h83db;
t_buf = 16'h9544;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2281;
e_buf = 16'h0000;
n_buf = 16'hcdff;
r_buf = 16'h3200;
t_buf = 16'hc2b6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfde;
e_buf = 16'h0000;
n_buf = 16'hd037;
r_buf = 16'h2fc8;
t_buf = 16'h713b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0359;
e_buf = 16'h0000;
n_buf = 16'h9643;
r_buf = 16'h69bc;
t_buf = 16'h99d4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h41c3;
e_buf = 16'h0000;
n_buf = 16'h5b56;
r_buf = 16'ha4a9;
t_buf = 16'h11f4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1f7a;
e_buf = 16'h0000;
n_buf = 16'hb9af;
r_buf = 16'h4650;
t_buf = 16'hefe9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9a43;
e_buf = 16'h0000;
n_buf = 16'h6a17;
r_buf = 16'h95e8;
t_buf = 16'hfb94;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h23fb;
e_buf = 16'h0000;
n_buf = 16'h9008;
r_buf = 16'h6ff7;
t_buf = 16'hc724;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc8bf;
e_buf = 16'h0000;
n_buf = 16'h5898;
r_buf = 16'ha767;
t_buf = 16'hfc15;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h69e2;
e_buf = 16'h0000;
n_buf = 16'hdba8;
r_buf = 16'h2457;
t_buf = 16'h088f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h27e9;
e_buf = 16'h0000;
n_buf = 16'h0067;
r_buf = 16'hff98;
t_buf = 16'h3c4a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h283c;
e_buf = 16'h0000;
n_buf = 16'hbf02;
r_buf = 16'h40fd;
t_buf = 16'haa15;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd7a3;
e_buf = 16'h0000;
n_buf = 16'h89d9;
r_buf = 16'h7626;
t_buf = 16'hb031;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h7a8c;
e_buf = 16'h0000;
n_buf = 16'h9ebe;
r_buf = 16'h6141;
t_buf = 16'ha21e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6106;
e_buf = 16'h0000;
n_buf = 16'h8a44;
r_buf = 16'h75bb;
t_buf = 16'hebaf;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h178e;
e_buf = 16'h0000;
n_buf = 16'h0129;
r_buf = 16'hfed6;
t_buf = 16'h5b17;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h953c;
e_buf = 16'h0000;
n_buf = 16'h9f9d;
r_buf = 16'h6062;
t_buf = 16'h26e9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha436;
e_buf = 16'h0000;
n_buf = 16'h6b43;
r_buf = 16'h94bc;
t_buf = 16'h46c0;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4b5c;
e_buf = 16'h0000;
n_buf = 16'hc954;
r_buf = 16'h36ab;
t_buf = 16'h578e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h79cc;
e_buf = 16'h0000;
n_buf = 16'haf4e;
r_buf = 16'h50b1;
t_buf = 16'h9120;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb7d7;
e_buf = 16'h0000;
n_buf = 16'h9cc9;
r_buf = 16'h6336;
t_buf = 16'h94fb;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdfcc;
e_buf = 16'h0000;
n_buf = 16'h6c9a;
r_buf = 16'h9365;
t_buf = 16'h516a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb4d4;
e_buf = 16'h0000;
n_buf = 16'h54c5;
r_buf = 16'hab3a;
t_buf = 16'hc95f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2e70;
e_buf = 16'h0000;
n_buf = 16'h1bc3;
r_buf = 16'he43c;
t_buf = 16'ha743;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hce9b;
e_buf = 16'h0000;
n_buf = 16'h7549;
r_buf = 16'h8ab6;
t_buf = 16'h5a43;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h30ef;
e_buf = 16'h0000;
n_buf = 16'h1c04;
r_buf = 16'he3fb;
t_buf = 16'h9a28;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h786e;
e_buf = 16'h0000;
n_buf = 16'h9990;
r_buf = 16'h666f;
t_buf = 16'h3a9a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he97d;
e_buf = 16'h0000;
n_buf = 16'h5e42;
r_buf = 16'ha1bd;
t_buf = 16'h3152;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h10fc;
e_buf = 16'h0000;
n_buf = 16'h0729;
r_buf = 16'hf8d6;
t_buf = 16'h4a11;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h3ff7;
e_buf = 16'h0000;
n_buf = 16'h4404;
r_buf = 16'hbbfb;
t_buf = 16'h626f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hccc9;
e_buf = 16'h0000;
n_buf = 16'hcdf8;
r_buf = 16'h3207;
t_buf = 16'h958f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2c21;
e_buf = 16'h0000;
n_buf = 16'h652c;
r_buf = 16'h9ad3;
t_buf = 16'hbbc4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h15ab;
e_buf = 16'h0000;
n_buf = 16'h3ac7;
r_buf = 16'hc538;
t_buf = 16'hd03f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2a7d;
e_buf = 16'h0000;
n_buf = 16'hae1f;
r_buf = 16'h51e0;
t_buf = 16'ha87c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h843b;
e_buf = 16'h0000;
n_buf = 16'ha2a7;
r_buf = 16'h5d58;
t_buf = 16'h7d90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hec4b;
e_buf = 16'h0000;
n_buf = 16'hb79b;
r_buf = 16'h4864;
t_buf = 16'hb1b9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hde6f;
e_buf = 16'h0000;
n_buf = 16'h2d5d;
r_buf = 16'hd2a2;
t_buf = 16'ha48b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h24b6;
e_buf = 16'h0000;
n_buf = 16'h5cd1;
r_buf = 16'ha32e;
t_buf = 16'he73a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hea5f;
e_buf = 16'h0000;
n_buf = 16'h8cfe;
r_buf = 16'h7301;
t_buf = 16'hde0a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h27f7;
e_buf = 16'h0000;
n_buf = 16'h3a51;
r_buf = 16'hc5ae;
t_buf = 16'h68a6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0a17;
e_buf = 16'h0000;
n_buf = 16'h959f;
r_buf = 16'h6a60;
t_buf = 16'h191b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9eee;
e_buf = 16'h0000;
n_buf = 16'hdc0e;
r_buf = 16'h23f1;
t_buf = 16'h6229;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h10fc;
e_buf = 16'h0000;
n_buf = 16'h2e47;
r_buf = 16'hd1b8;
t_buf = 16'h1b9e;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8a8f;
e_buf = 16'h0000;
n_buf = 16'h13ab;
r_buf = 16'hec54;
t_buf = 16'h1b92;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h399f;
e_buf = 16'h0000;
n_buf = 16'hdc6b;
r_buf = 16'h2394;
t_buf = 16'h1c90;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h1081;
e_buf = 16'h0000;
n_buf = 16'h308c;
r_buf = 16'hcf73;
t_buf = 16'h28b4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2168;
e_buf = 16'h0000;
n_buf = 16'h1773;
r_buf = 16'he88c;
t_buf = 16'h17f3;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdc4e;
e_buf = 16'h0000;
n_buf = 16'h7e97;
r_buf = 16'h8168;
t_buf = 16'hfa69;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0a66;
e_buf = 16'h0000;
n_buf = 16'hcc66;
r_buf = 16'h3399;
t_buf = 16'hc788;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2df0;
e_buf = 16'h0000;
n_buf = 16'h3ed3;
r_buf = 16'hc12c;
t_buf = 16'hcd53;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h4cea;
e_buf = 16'h0000;
n_buf = 16'h8d10;
r_buf = 16'h72ef;
t_buf = 16'h6482;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hba02;
e_buf = 16'h0000;
n_buf = 16'h95ee;
r_buf = 16'h6a11;
t_buf = 16'hcd0d;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h03e9;
e_buf = 16'h0000;
n_buf = 16'hcc0e;
r_buf = 16'h33f1;
t_buf = 16'h84ee;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2fd6;
e_buf = 16'h0000;
n_buf = 16'h17e3;
r_buf = 16'he81c;
t_buf = 16'ha5e6;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hc247;
e_buf = 16'h0000;
n_buf = 16'hd9ed;
r_buf = 16'h2612;
t_buf = 16'h1b98;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h6a1c;
e_buf = 16'h0000;
n_buf = 16'h0a15;
r_buf = 16'hf5ea;
t_buf = 16'h588c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd80d;
e_buf = 16'h0000;
n_buf = 16'hd102;
r_buf = 16'h2efd;
t_buf = 16'hd58c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbc20;
e_buf = 16'h0000;
n_buf = 16'hbdb6;
r_buf = 16'h4249;
t_buf = 16'hcb70;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h72d6;
e_buf = 16'h0000;
n_buf = 16'hee52;
r_buf = 16'h11ad;
t_buf = 16'h6748;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd505;
e_buf = 16'h0000;
n_buf = 16'hf341;
r_buf = 16'h0cbe;
t_buf = 16'h394a;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h54a1;
e_buf = 16'h0000;
n_buf = 16'h415a;
r_buf = 16'hbea5;
t_buf = 16'h2a7c;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hb353;
e_buf = 16'h0000;
n_buf = 16'h3dd6;
r_buf = 16'hc229;
t_buf = 16'hae09;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdca5;
e_buf = 16'h0000;
n_buf = 16'h084f;
r_buf = 16'hf7b0;
t_buf = 16'h9518;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfbd8;
e_buf = 16'h0000;
n_buf = 16'h96c0;
r_buf = 16'h693f;
t_buf = 16'hb8ef;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2922;
e_buf = 16'h0000;
n_buf = 16'hd77c;
r_buf = 16'h2883;
t_buf = 16'h0a12;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h19ab;
e_buf = 16'h0000;
n_buf = 16'hd1ee;
r_buf = 16'h2e11;
t_buf = 16'hb144;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hccf7;
e_buf = 16'h0000;
n_buf = 16'hf18d;
r_buf = 16'h0e72;
t_buf = 16'h3ef4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h08b9;
e_buf = 16'h0000;
n_buf = 16'h2b01;
r_buf = 16'hd4fe;
t_buf = 16'h5da4;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2619;
e_buf = 16'h0000;
n_buf = 16'hac51;
r_buf = 16'h53ae;
t_buf = 16'h3ca9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hd43f;
e_buf = 16'h0000;
n_buf = 16'h3d26;
r_buf = 16'hc2d9;
t_buf = 16'h37fa;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hde62;
e_buf = 16'h0000;
n_buf = 16'h1209;
r_buf = 16'hedf6;
t_buf = 16'h6e66;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h195c;
e_buf = 16'h0000;
n_buf = 16'hd512;
r_buf = 16'h2aed;
t_buf = 16'h64a8;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha7f5;
e_buf = 16'h0000;
n_buf = 16'h154e;
r_buf = 16'heab1;
t_buf = 16'h22a9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hbc20;
e_buf = 16'h0000;
n_buf = 16'h5db5;
r_buf = 16'ha24a;
t_buf = 16'h9179;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h75f2;
e_buf = 16'h0000;
n_buf = 16'hde3a;
r_buf = 16'h21c5;
t_buf = 16'h07c9;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h0e7f;
e_buf = 16'h0000;
n_buf = 16'hd656;
r_buf = 16'h29a9;
t_buf = 16'h295f;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf7f6;
e_buf = 16'h0000;
n_buf = 16'h0445;
r_buf = 16'hfbba;
t_buf = 16'hf135;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hf320;
e_buf = 16'h0000;
n_buf = 16'hba8e;
r_buf = 16'h4571;
t_buf = 16'h6470;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h5f0e;
e_buf = 16'h0000;
n_buf = 16'h73f7;
r_buf = 16'h8c08;
t_buf = 16'hf206;
nprime0_buf = 16'h0000;
#10
m_buf = 16'ha8f4;
e_buf = 16'h0000;
n_buf = 16'h33db;
r_buf = 16'hcc24;
t_buf = 16'ha4fd;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h8147;
e_buf = 16'h0000;
n_buf = 16'h03ba;
r_buf = 16'hfc45;
t_buf = 16'hd8ed;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hfe39;
e_buf = 16'h0000;
n_buf = 16'haa40;
r_buf = 16'h55bf;
t_buf = 16'h062b;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h61d9;
e_buf = 16'h0000;
n_buf = 16'hc10f;
r_buf = 16'h3ef0;
t_buf = 16'h9d89;
nprime0_buf = 16'h0000;
#10
m_buf = 16'hdd9e;
e_buf = 16'h0000;
n_buf = 16'h2284;
r_buf = 16'hdd7b;
t_buf = 16'h8f40;
nprime0_buf = 16'h0000;
#10
m_buf = 16'he6ad;
e_buf = 16'h0000;
n_buf = 16'hc16e;
r_buf = 16'h3e91;
t_buf = 16'hd5f5;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h798f;
e_buf = 16'h0000;
n_buf = 16'h816a;
r_buf = 16'h7e95;
t_buf = 16'h23da;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h87a1;
e_buf = 16'h0000;
n_buf = 16'h47fc;
r_buf = 16'hb803;
t_buf = 16'h7185;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h2923;
e_buf = 16'h0000;
n_buf = 16'h1d03;
r_buf = 16'he2fc;
t_buf = 16'hfa46;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h809f;
e_buf = 16'h0000;
n_buf = 16'h3fe3;
r_buf = 16'hc01c;
t_buf = 16'had98;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h9850;
e_buf = 16'h0000;
n_buf = 16'hb476;
r_buf = 16'h4b89;
t_buf = 16'h1965;
nprime0_buf = 16'h0000;
#10
m_buf = 16'h044d;
e_buf = 16'h0000;
n_buf = 16'h84c5;
r_buf = 16'h7b3a;
t_buf = 16'h149c;
nprime0_buf = 16'h0000;


	#100
	startCompute = 1;
	#10
	startCompute = 0;


#10000000
getResult = 1;
#10
getResult = 0;

	end
	
	always begin
		#5 clk = ~clk;
	end
	
endmodule
